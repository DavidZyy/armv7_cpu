/*
  control and decode unit.
  decode the instructions, and issue control signals during
  different cpu states when executing an instruction.
*/
module control_unit (
    input      clk,
    input      RST,
    
);
    
endmodule //control_unit
